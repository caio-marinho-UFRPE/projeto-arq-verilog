// Grupo composto pelos alunos Gabriel Leal de Queiroz e Caio Vinicius Marinho
// Atividade da segunda VA de 2025.2 de Arquitetura e Organização de Computadores
// Implementação do NÚCLEO MIPS (TOP-LEVEL)

module mips_core (
    
    

);

endmodule